module rob_testbench (
);